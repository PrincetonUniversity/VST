(* Copyright 2012-2015 by Adam Petcher.				*
 * Use of this source code is governed by the license described	*
 * in the LICENSE file at the root of the source tree.		*)
(* A top-level module that exports all of the common components of the framework. *)

Require Export fcf.DistRules.
Require Export fcf.Comp.
Require Export Arith.
Require Export fcf.Fold.
Require Export fcf.Rat.
Require Export fcf.DistSem.
Require Export fcf.StdNat.
Require Export fcf.DistTacs.


Open Scope comp_scope.
Open Scope rat_scope.