(* A top-level module that exports all of the common components of the framework. *)

Require Export DistRules.
Require Export Comp.
Require Export Arith.
Require Export Fold.
Require Export Rat.
Require Export DistSem.
Require Export StdNat.
Require Export DistTacs.


Open Scope comp_scope.
Open Scope rat_scope.